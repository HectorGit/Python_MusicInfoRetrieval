BZh91AY&SY��7L ��_�ry���gߴ����`S_  �T�UM�� ����C@УZ��v]4�4m�ff�1��];w6mu��f��҉�!k��if���f̪Jٶjih.�mTP�6�&�P��Rr��J�"�R��6,
֕-�8Н�`U�X�p��+fJ���kN9����cm� H     �~���T��0�i�!���M1$��d � &� �����(ڙ3S�f�F@m ������j�J� �   � �&M4�dd�т0�F� I��A@��2&&�M=!���zz���÷�˿˪@@�<�B
@�'Bd'����@F��~����ʏ��\�f����$��I �s?TR�O�$�H��l�h#,Hp���4GD�V$�C�>�G��}w�+��}ܸ$20	��Ca 0�X���!,`B� X�%� X��X�B�B 	c2�$��X�B�0�bBKb,a�B�	b(HB�HK��!b P��JX�IbBK�,H�P�Ig�Dm������΂�|7>2��iIێ_N�Bg:[V��o�?�g���+=5Q%�Ȫ�ڕ*"v�N֊wX��fU��ܺmhu�4Ӕ�����U(RV��ɱVT�GdW����[&C��;"]�����w�����q80�u��yUx�`���ד�&Η�v!r�n��cfŃ���aM�e6���K��t+jk��E�Ж�v�j-�yu
��ބD����Z�impڅ!i\���mSn!��J����-��s�K�śV ;O\Vv�-��*����3,�v���%4`�VjRd��2̫�;���J��{mU�KN�WF�;4�6ε�4�8L���R��,�D�u&f��9��Ԩ�z�k�v�~��s4dyH�ۘƢ�� �b���Zad*�=�d˲��+0n���sEGv��pX�(,,bVP![�(��(��b�9�h�6%��1T�]�Q��aJ ���x�4Yc-�ڷnb�=��N��D�0�Υ8�Ub�Sb�5��K��Yl^-c���cS*$�+���u
i�W�P����F�u\z�6�C(L��%3)xT�TF�B[��0"l�)Zie��6�ku1q:�w�Ź�YD�ar��b��UĦ�fQL�e�(iyo�!ie�S7�\�Ե��Z�DXĈM��� -ΛnF�֦�V����<���f*��qd��2Ф�pk��Vb(��Z]�I�h�1i8�*�Bl��[��
G����LV�]ͼ˦2��4��X�5�f�ǻ��]ч3)���HƩ��&-��dd��6�,�Ys0������˫-ۼ��(�����#�$�$��'�R�Sqp�i9��X3R�W���`���r��Y�.:T�2�w��;�q�e%[s����+��i�.l�na�ɶM�2�����tv^b����Z7�SVݷ�*��
���N�*�˒�6�$��Y�rPÒ��[a}}lR#�Yq��P��x�/4�N}X�䑗K�����}�-ٲ�k�����n�z��k\��#����O�<�ߞ:ګ�[?D]�0�y���g)"��H`�W�X�����;4�wC]��1b	�:�o��a+��'d)�qZhTm�LLeH$��j
��t��:C�`��r��h���ù7\��[�awc���r5�r����+����v��5���6����{)-0_j<tV:Ҁ��WX��nt���#2�1ǁGs��� ޣ-�ަ�Gd��Ǖ{�hk���f��glƁ�'j�C��s(�p��*�\kr�k#)��xl9��;�[�Nt�4f�ǀ�](�ڳp��+�:�K�+�[��m��f��م��+z��r�^!��.]9�5	����G�]q�&�b�|L)ηή�,XO\|��[�S���o�\�;�%p�&*w�������aV��1-iX�����v9��b�W$�':����?;�=@��7���R !���/cU����>Ԗ��&�ڍ��FfZꭶjwS����K�՛�_�i*�MJ�e�K�c^�������({S���ĖUb��U��1_+�޼����d���t�L�]8�reZL���i�rX�J��k9К0����rb�����HX�*r��������CTEc�h�;]C���m,�*�5�f�3�k�E]�L���+D���R�=J��PW��Sݕ8���y4i��Q�$�oI��/j�(�cYOd�ț��B�����kG"�;�m����7.�'�
 �]�j��,`�W�f"I���u�Sc]{��λ�v����㽧�"��県��zd/F9�'w����;�6vm�B��2C�?1�0^�t.��0<�8�v+x�p�*fdس�-��Գq�N��td�o�B�x��b���r�s��u\qg(.�:o��=�vp�ӳ��+*Rm=⫅�
��[&�La2d���{I�ɺ�N�5�$�I,�ߝ���Wy�� ���8�Қ��-��&�?��j���٧�$ 8��َ��]{ �9m���^@!�9�Q�&$� ��P�����>�N��?��5���^D2��u��B���'����w�ߔ��-.Ӏ�{�ѵ����HG���0vt�wV����+]
�Q���ș��	%�+_���ɩ�&L��uuuuZ�\�T�K��E����a��J�v~�{R	�v7Osw*d��}�!�.��\I��i{��;7��@�I�#Ӕ�Y[��Ǝ�-�3 ͎�|�W�N�ut�*T�N�����uuu*]Rm�9�S% �	a�$v��˛�ù�̬������e[Ⱥf:��)�.�J�-@C.bL,LfE��5�"����F˕�A.[��}�����]]J���������6&���j��n��c%ކ+�e��y�z��۟����+Qg1Z������#c�U۳M�HO�u1d�]u����cb%���׋���Z{3���vL�@Њ%���4CK��L��N%fZ�sv��kkVK����v�����l���<��sa�UrVTv7,u��]t�a��J��n.XF(�)�4�UⴜI����;��Xk�`6i���u�R	���E|�ڊ����L�v,�[����j�.�q���9���IS�^���7���!]�}Z��Rf��D�U���/�HQ͗v�� g)��p�2Ƞ�x�S��0nPc��/)+٧��+m��Wu�u�'VQ��7`���	L]�	�6�F��w���w��}�D|��u!��G�×���BT�qr�"�)�� 0�P��wy=�U�v��VJ�XVfg�Q4K@u�#�a��ʾA�l��m�<���۰��[Ө��]�':ċ��y�/(wqO�(V���:�������C\4������6�'��S�e��6-嘍=coK�NݘpKNq���x�'vt��	dG�]�sj��FT�K���s8v���1�t���M]��Wl��B�p�e@R�ƻ\jr�G��sWסLb�wN"����x��v%�u�MWӫ�~ U�%k�T]�ʾ�A�z����UUI  �G��d�&��Ma�fj�t�����9�_e�f����o��K��dy���SK'@і�7��v��<եY��|L\N�O ��0�+k(h���;�w�H�n�Yq���o䎳
V]�t�a�̌矅��w��rT�
(�d�A��PXh�UQH�X��)UX;U���QH��h=�6�^�g4��r��+��}����*�&v>��*hX�}����E u��{2����ޙ��ޕ��z�ǉ:��u0.^��unz��X.KdLg]��o�@��Gή
5�8x5���B��8ʼ���k$C�i��b��+"1�*g���M�V���S�����Lg�];�jt�Y���S��U�wKS�:�X5�0�2N7s�x*�?OoT�^�Bn~���8�?��CF4Y�e˞z�c���k�<��k�ە6a7��ր~՞��S�mz���u�����n'��L�@U]�s@c�'X��٩�6�p���ȧo9��
��y�4�A%tsL(�ڼ��u�p���_X6�=͚�*9z}X6Ա�Mj�(��~L���7pˏJ�$�i��*��xgg����YR*`�[}�x�[���贇���c�}�ez�ޮu�+q`j���!�`�:f�e����(���TO�jI����G��޾�(�<&rt[�]CE�+=y��]<�zA�մ�c��(�f��-�B���������/�Ox�6���N�ꀥ[��.]���R"� �D�#�߮��EG�H���2�!�Tj<���A�u���s�J��]���u���m�m��7�>�.�v�?z~��]Q3E=���*��c�\�yQN�i�Kp��ҍ=D΃&���¡{�4�34�������G�����"b��fp~�i���dcՆ�S�[��S�����rEu�GRv�v�/,�T����<��6�]Xޭ���Ru���\��m��e�*�2R��5ĩ��ݩբʠ�!����'aw[�ʹ7��t�Mn��i��.i\�m)[�ӧ�C�`$�%�f��Ԯμ�}O���2V�;]w�ۀ6��!���/����Z��7{��4,�0#)��ɓ%�	��#��XdA�D��#J!LR)�Ib�b1��?Ө��SBs�c��#b1�� Q��|G�ǂ��N�So�ZD��R��.56O�\�Dϯe����Q_w�i�X���MJ���aW8�����eZ϶�ŧsl(�-k6�jJ3+�X�B����^(��/��#��\�d��j�i�O�������l�F�h
�Š	�*�s��i���P�c��X���<��z�~>o��)���<ױ��B�o;�����E0���z�8�~a�۲�����z�ˇ���|2�A,�0���~����5-��B��C��aء��a�3�Z�W0uHr��Ʒϊ�籯=����~�U���R��.���b,ə�n��5���[X�
v�>�OR-/p�g���{��>2��e)�����i�\�o{5̜�DA� ����{h���.��!�'�|v���5�9/�� ޯ�X��;�ݪ�s�#���[9�F��Us�XH�W&��.'��a����*v�o~8j���H#��ff��GE���?lq������btUՌ(F]r9&Xb3`�N�~��c��E`�_�8��썻Y=�~/���,Iz���o����Śs!�dB����7��+?D?Y1ƿ]x�����Ժ�ۄe5����SI��g Tg���b���jE�fs��F�>��!9^��ܗW;dsP�}�7�y�{���dP�o1�z>Vfn8%�k'��C�����s�k����V򣋦�.�}-�lj3x~�[Y��z+4���L�����33E��#91鯀y����c���Ϙ[0e�}y�/��5�����v�h��b����s�:$��>�c'�n���:�N�ʠ.�)%��37�3�h�\<`���C�ʏ��O��gR��C?�pe����U3Y|��{�5b,d$a�������DDB�n=��,�O 3rH��7 �Q�� �Ӈ���rnF�mf9e�� ����fL\1t���B�� &Hw���ՔI͝�I^~2�M�ň��]�|���8Q�VcW��ء�,��#�1�.����?L�2~�1��~��%��gf�V]���D2ւ0��ެ�݂ɴ��Iv��&=g�2U�۷�)�+w�
f�Ah5[jgw6������r9��6�X�fJ�EDP�ʅ���q"�i�Z(��D[LQj�QD���ƪ��B���UV���[�Ea�BҚ�N\�sls�ֻ�5OB4���?W���	�i��N�J�]��tf�p�i��dǀ��Ǵ��� �z�Ѧ�n�K_�\��\X��U�u�(�Yș9hbi�o}��}�GO�g��h�?\U*TK�H��N�E�+;��M乭��X٧S/-�P�1�����0��t�q�9g25�6��n�n�ɮ�yɦJAK����}����.��֒���x�O��f%i'i�l)�(�����F7�B����ә[Ǳ���k��y��h��-B���c�?fg�RmQ~4}[d{�b3��{Zjs4�2�B7D��|!�=�'n@�T��G��י7^|aݏ�cc���Ԕ\�Pŉ����*���@�����HW�mq1��� I�d5z>ΰ����;:2� �9+)a�$)��B޵)�>3�(C�Z|<=i�k�u[��}�>�t��s��L��ffo���yE�L��̀*�9�W�*�mө�w���i/^g�!�j�g���y�tq'���㿚N�W�o����S�N&�ȅ�;������z�n�EO)/1dx�8�{��^t�F�E]*'�e܎7��~�> Iud{��UT�Ř�S���s��Z��&7T�Xۭ!���37�U-���!��|]����e�e�jW׆�����K��&���gWyM�8�c�ׁS&���d�i �;τdM�3U��]|L	�3G�T.�3���7������P��Y�Y�߱�1W��gk���������r�iW$d0KsL,�fTo��=L.�~��V��\�;띵��M�y��2�t��grk��C���X Щ�fy��p�u����;�Z�1�5��y{��\c�r���;T���d#j���������uޖYv;AF���Ba�������<)d�F]�[u}�v*�V	ƈ���B��uT��DcP�iV��aL���Bv���;K����c�G,�����v��ΧM���{����aŁ;�}g��k\4X�12����9:��	�D�Nd�*�D
٘���(p�D;�I˽��męwZ��9�S���,���/��0��W�]���)��c�R��KTAqTa(UpQm�SQX�ݚh`����4�.���*6�UwAH���`��w��f�Ԫ�M(�,cZE�"ڌ]�Ӗ��]4�F^�:r��G�{?*�^�M��=�f���H����b���Ҙ�4y�d�8�'���}Y(myv|�!ӟ,0;B{��f��7.X��&�������߻BFz�\��d�,��gC���/�%V���}W��P�3��W��Vƶ^*9 l�x>�,M��.4}x<=*��߾a��h�=X�r��f��=���'�s���ns2��4;�hؖyژͻ��cb�-�9um��߲	�p�4~}���~�y�*|����YA��CN�H��0N[�o:@��G����oY�/�6��;i��W�04�U�TK�/UoZז�		�nؗ�9Iy��N�5�Ϻ�޾����A(۵�[s�W�zy�����}F�F~���S�Y�!��LZ��5#G����a7&��l�M���1��g�,J�:�hQ�&���~TfWizP�6,g��4e�_����j������'��]uC�Bx���g�ީ��H��M�ɣfg���9��75iЛ�Q� \Tܼ�b����14���X��Q3�6�b� U�z}mf��G��t�^ Q��S�o�ֻ�����|��Vp:��&I����}��Aʎ1;M�L�+1��M&�t�0?���t;�o]i��h�(���׆0�JA=��g���"h� �T�5.;#7T�_wE�1�Z��AQ��}�.�`sM���@.:\����L��{^���5WN��+���� ��C=odRY3P�Nۙ4<U���}���|�/\K
��M�ބ���Q���zb��uE�͝�H���~�o�L�r����M*�7-(\!�s����5tܝ�߯��^�9ʫ�e�{�
�/H������XQ0#��s5��qȜ��s2�c��5Ār@/	��S3@�W�)�s��5˛��3]F9��v�mb�.f�),R�qnf V����2X��m���hѮ����u/f�#�ie�	"m&�4I��vU���Xuw�. ��Уo�I�_�r��T3�w�R��ܴ�P9S�GF[y��]�Kmr
����K=�Ո)]YtK�份帅VJ��-M�3�]�a��0n`ϻIUR*�E�*�B���Yn-��F�b˱��hT��Q%RUP%P�FR�,JB�"�6�-���wv�R�j���.(��H���J��rh���0�`LLǚ�G����o��h���r$�<vU��)�f��6vb��m�0�;�!X7QەVG��tՙ���˾ʊ�_���2&V��рX")'��|��;�.L�����M��"�{1฿a�H�K�{٘F��4�L��(���/0���X�P6h���8O{j�s��4�W�'i�B.��������t��P|�������Im����=(��u;gԦ�m�T{��ma۫ q�׬�3,�>�YA��%>����&���u�Q��*���đ�苾�^7^�ji�V#��{t0�6��[ؙ�FK~�.$r��R���&�TY$1^b�TP��>�t	��{�P8����V	I��̈́�d~6{�<���N�G�q	�'���b���X��+�30�X�E"r��M�X�%u� ��)6�O~�]L��g�'G���X��W틅�Etb���ސ�RX ���ܱ����ʎ9T��~o�2�������B|a.:��G�'�m��b>���´#���T�68Tk!3���)�x1N��=u�����U�M�h����e�]x'gW?_y箂i�dɮ��].%פ[q��j�@��0�Z��"��E�U�a^�_����[B�?��,��Tݴ�֤������wbsΩ�f'Z��g��bO��0��?QՍ������;�ȸ�W"��&����y�;[���s}B̛���Q��1��yq5��2���e���x4|����gE]V��V@����J�?z}�Q�k��QJb�0?H�U��t��[2���hC=�O���1�+*���ަ����{�����Ҭ���,�砒����j�����=���Ϸ��K��8Q�E��y��_l`�v'7aíșf�SH�	C�S�E$阙�L��h.6K���e_n�9n�Z�/;�S��Pĳ�����2�i�˭��k:J�N$a;0S|#�]����]e>kgB�tW���1�^��E%_%�0�ݭ��Ql���k��͊��%g?s�+������M,:��ﳦ!�S�/��B�]e]��R�P�B�QQ�������V����(�J����T����KZYWTR)Pb*�QAEZ���SO���8��ڻ��c^�=�?�v�=�5��w�i�t�4^zج��so�J]�:��y=�<N��tg�s��������U�y-u8&�нr6?���zN/�J��Q�?��6i`�j���LT��?���;��mz}]u5o���)� `|�48���ū4�ټl�"�SSڪٞ�p�n̆�D�o��D��C[��>��yn�M�.uFzz:}ԞO��/yi?u�`��=��E�x��5ux�������`�nZ�0���Q�ŋZ�����ټO����x���b�P�rix��u��0ve^\��.O�ty{8<DI,�M^>:i��}g���݁�z����4�4�Il7[e�sF��cd�|��%*{f~�p�����^�R5)_�S�V]������]K������U]&Q��S�kv+6-�`��l�������5�]?"i� ���O���]u�e��6�P�]d�9�q�iH�`�^oR���H{��$��g�W�RQ�9�"�&�z;2{yu�.���ݼ��~��PΙYY��E��6�(���,T�9���D��)O�sa#�gz��{�4�P�n����3��d+��x��f��f,�L\�&��5��ix��&Nh�fK�\��e[0z��-���1L��`�껡��
jګ�9O4�u3�0BN�}Z��������N�X��g�fW���f����8uP���X�똄A�.dB���Δ��'G����yx��ȟ+�k��3���To�*���j�XN^N{G������������2K�0	�����(Wr�t>���PQ��ڀQõx��V�PCjܳ���Y�4��2:u�s^RL�3R�\k:��Z%����c��v�噻C��pNo{�1��V<(�`�s��ظ�%R3Ws�B;VsY��:|]]բ45�u��̾ï�,��xc5��3^�;`���U9l#]�%�ޣ���ǭ]��'�zbO��TQ�W��QFDQh��db ��F"�`"�e�4�ƚ(�
(�*R�B�9��(c�Q�� �JhTxw���M|����GMx����2����N<]�����W�u��W�G��N����gn��u���ʯ�$��a���������ʒ�^����{�^!'U�j�/��y����j�Y��U��W6'V[w9P��\.뗤���~��RH���n��C�N���a�>6s���NV�=2��Eg-�Ev�����w�������v�vE}��֊j4��������КUs�<'y~9G*��*t<����	�{�i?}Ɖ�^��MG|��O�H��}h��v4�6sܝ�M�T��&;�I����+�����u5�MB����7�sN+.��a����c��]o��M�O�0�.&�f�$�<Sbax���c�R��$�y�.ɂW�~6��E����}S�l����������*е*+�wK���Uv��ͽ[s9	��B��_�鯫b)�}U8�2�"wb��'�f�.�Q�i�є����[d@W�$��=a̔.�	K7�uIjt���YO*xT{�u�"gس�Xp)-uO�b|>�G��ɒ��;��1{��/1��z�0���6��f�W�+�}�������^��<�%���)��|�n���Yw��9��ܗ�j��*�M��0[���5y+�^
	[پ#��m�ؒ��]י�-�u-rվ�UM
�~�1�zX�#c��*'���fƔ�`��R�2�=⭫�X㣕<&���:ؗ�@z8��]}*�c���qI
���}��W�(�n��Yz��Og:�Pw��Lٺ ��X�f�fɘ�����0k�D��ݪ�(�@�����5&�R��	y�l}�N�d"dls�@���l�JvF�5em�B������� �!�J���c���A+W�:�k�$XI����/T�	C���n�M#�M���)��*|����&����!Q7	F47N�)؝�%1i���n9�z�.\sOI^$�>��rl�e=���V7�Z��vΘѱ�sg8-Ъ"�1�*"�b�0�bb�b���b��H�D)-�ԩH��C��UciR�]��2m����$6���1=�ˋ�P�S3<u�:m�4����1K�8[���0����_�X��#��G��W��T��B&/�e])X�>Ǥ�+x�׶�槢n�Z����ήvF���ⷉ	]̭�I��M�ʐ��c�l�Ɨ�O޻�q/���Q�}�yOv	1��j�A��)O3��J���'�q�4Y��-]C�=b�fkl��
��������-�=6rW����������=����0gy��1j�E��5�w�h$���I�09<կ�Ԩ��S9�n'��#�)R#�g�Ge��<^�%�u���T+��糳�Vn  �j<J�Oj��;6��n�n�-��;w�����pǲ`��a��ή���33�	E�����,�M?sŒ���Q��[<U|x�K{��P{=�]�&O��V�l$bX��,��um�'?Z4P���[^�̨@��0o�!s�7�c�#�j���}�@��J��7�;��zu]�d�݁�+b��QU� ��@����ƛ'�����R)R�(w(G/8�`S.]�>u3B��\�Ȅ2���uX��p8��OZc(ʃs)�������7�<�_�*��v6��1��P���D�:X!��:���^��\��DƱ�Ø�S�~�Jlک�+�:�(���
�ۚY}��E�� ֗1ˮv���n�0�?��幼�nk�������J��4"�U�筊�W\�t�]��Ӊh�)�Lj�գ��>�ɏ%=a�d�,�V���ꏗ��
h�r��|�F�XP�q�F-��*kK�w���k�k��κxj��X/~�f������u���Y7��u<��w��U��*g�5=#Uk7c:N�j<�v�Gwݣ��(�p�e�j�6�dꐶ��y�e�@Ɍb
��7�k!�Y������yV����>�e��8����L�;��N��{w�xv�x��"\�."�i���v�a�����cλ;9\sv �����n2Y��*�<9\\o���۞�J��B*��M�E(�w
JTUQEU��Ub�PDPDJ����������QV �TU�k|�c�b��3�3uG�~F^�?���ʔ��p�Wj���]G�5u榩|��W��j�x����Pvb���<C�n�~a���I���U#Hx"W����ߚ-��^�7� b����L��ܿY��;1p[�q��e�k�h�\���
��MD�nen��Նq��.�cN���	���/�\"BƩYO�
��p�Ԇ[6p{�z��A.���P���]�\f��mM8�}���&)Ʋj���Jc��"�@���h�u�t]sN�
N�+��`Z+�)��T��
v׿O�r�}�`�j��o�T7�\?v-�~cL:�����L%�w�N_&��_�ɘ{2�a����e�z��H�G��yR�@ͤ�;id
O��'�U��	-�PR�ٞ�QQ/ۣ��
ҡ����gͤ���Yȫ�d�l5P̺�^G=V��S��p'���>���zu���!H��QHUB��6��L$W�螆}�E��3;{T�(O�&��������z����ux�Ԥ��p���/-��%+Q�聝�ј�b�"�|)m=!T�b��U�������6�KH� �SC��|�~��s�޶��(�؀]�ɠ��{��>^�9n�##6ұE C{3�f:��!/��p��U���vG}7�"+��t�r��8k����瘬��4V��rߎbu|��:q����H��]FX)d`�u��9��(��Mς�ժv�̉�h�{ۧ���} WO��3
�`���3C*�Ǡ>_z)�4&��h{��C��c��9�zNUK\��qH���hT���	��h62 %`�sL]{躓g՗�'�L�^��MC��0�f���]FƖV]4�ʫjb�i��QV���Z9Ќ���"��~���Y�)w�DF�� �L?��y��_�ڍ�E��͞�l�0�-ul�:J޵^:i�jd�"�F����tl跂Ĭ�xB*L�e��]�ѝ+�yM(���@j����z�=�\쪺��yU�
(]E���.�UDb�RTR��Q`��$U����u�GSv�D�H�Z��L�����2ݳ����6	�����p^���ݗܷ\Y �qZ-�r��@��T�l�.�����t"���B�-�h�elm�S���V�x�k(g�̻n����|��/���R�dt��.)�l
uR���B��"�������B�li�h��պ4Mk��cL�z��Њ���W�����[֮�Գv_�5\'�=1�2"���'ў/�,�Xˈ&z�t�A5U]s���e�G�%K&�%�[}�|�^�a���9�r}-:}��ӽo[:i����!ۂO�/1!�-���W8�/b���1r���#�YǞ=t�\���HO�V���5 �N?M9���[�����C;Z�B�
�fӘ�l��i4R��S�S��,��.��
h3��	�.'�u�З;�`V.��7ܚ��V��"���M:�ƎTux9����?X�:�\�����)k�xy!:��o�%��)y	��uo���Ӂ@YH��1~Δ$׆ו<]���j�w�' �HN�-�~�8z�U�'�I1S��F������ʼ��r,檇R�w~�;1J��5�9DM��!e�~Y����݄�K�)�Ʉ�t�#c�0�.Uǒ�GF���񀺲6���b�G��s���<�)�.SN(���K�hǮ�R������sj�Wn��t���{�gA�F<��������&2L�I���=�sKV��m\�t�Q�0�'�$��@%EV�BI �����ݿ�a!  ?��qʱ\��`+ZԴv�K?k���Œ̉Da%J��D�C�!.�D##$�D�# ���X�%c%MY!hB��L$!�`�! L�B ]�,��!$�@�!%�$ ��A	%��*H��M�>��BL3M(6BiZ��~�����I�BHA@$A@�H�J�ʪo�J/�7G� �в�D�5k_\-}60��-&� ��Y#M�xX(h��Y��F%��?^�|��0�僿??���_�^���γ��I ?87�y��W���'���u�B |����Dd$��IH�*K;���:��Cƃ���d&��;rIrD�Ǘ�Q<Q�}�H�����I�w��E��X��Y	��e�Fͤ�0;��v����R��육��d�WV�i�N[_y�ò|�<����ĳR�$ /����W���EH(,�� XE PQA@X��"� ����
I00
B,�$�R��d*$�a He�
@��4dQYV2JF�zW�=?���W\,���B@ �%D�(DH"#\�И�(:��!*�������C�����8`9�� f�@�c������g�����QՀeHI C0����q><�`k?��������B��Y�Q8�d�����o�y��SìO����<u��K�'���o*�����pv�	$ �D=�{}�!c�hkښ��8��`#:Q��ډ �!$���O�n�|W�at&��1Y:J��@NF|���p�$̮�0��X+�I�F�h,	 ��jM
Cð*I���>9:U-QI?����$<2!��[�T.0��3LR!�}�!$��`�=�����}���zT�� '�X�v��b�� 9�� �{$�����]'C�ñB�Ǡ���y��C�s��B~8�{9��M�
��@��:�<O7�$_��9@��y�N���\�� T��̽f�9�Ǘ�&�6�@��y�h��1"N��Y貆"L�GE���wz��|{`q~�|z@�=x�.&���޽^}gI���{��i&?ﯱ�	$ �x����c�TQEOL��xc
�����k��ܔ&��Ć}&�)�GY�(�ڻ�D�t>�3 v�t�#  }�����7:�z�'�����7�t��ڳ� xG��0�Gu�nȰ�N%Hi��ʯQ���>f�$���ʐ=��@��O�rE8P���7L