BZh91AY&SYe�G �_�Px��G߰?���P�ǅ���
L���I�� i��4CSM  � h4  	��S�di�i����@ �� $�A�4      	"I�����Б��DL!�	x!�"��HA4I8����)0i-�C iy�N)!ne��^���6�~[w����>�x&S��+0�a�#�g.���ݕ��y�q6�0�آۊ%���Xw��0,���Sl�Fl^\\�"P��A�Wta���%
8�Q/2�w��d|��1��E�H�(C�R�G������C���i�7:���U��R�Vy�;�(ɘ'3X�P`s�@el޵PD�T�.V�ʸ�`�(@�Iɑ�����Y즪��l �$	��0�+\3=Y	�8 2���Rg�lEM����f�	/7�u��S+;F��'QZjȈњi�q�;^L��0a��5Z.�n�)�-B����"��M�����M�>�� '!�2 ��B [�AV����L���*A�hfWxtI�~�����P�8Td,�Q1��=hҕ>��ʾu��Q��/?��dK�{����>�� 4غ��oYo��(>�F�!A ����q�٨�4w��ھ�`�<�D��m2X����� ���Y�M$���x�����e�ɤq�o�a�V�6@��a�8�ƣ,���f��`y���4,j����Fw��NE��`Ud�"�fs1R3;_#v	��Ex�["�d���QI@�D�\�4ĖV���K�q�����u�^Ɇ���v��TL�e��7��!�Y�X�a�P���h�J��Lh0ÑpcEX��(�fl$d�B(F�%'oO�NR�cX�&�1��2b,#�Ȉ.�;KA�<}>A�d{F�@]��plm8zĻg#x��"�N��u�;�&ÕX��s &9��5&��zVq7�+��Q/��7#p	�"Ku�X���6��9+��"���-X�DȈ&�(d:05c��5��0
Q�Q�>�cG���W�]��BA�
1