BZh91AY&SY�� �_�Rxg����������`�7��ܘ���g@eAv��5?H�6��L4�14� 4��Q=M4d  4  4 i���i��4�0LL��!!�&��='�=M�2244� z@�ᦙ�&�`L#��i���
�@� @4A�S��?T�i����=#OSv�BUJ;RL��D��!����?����G��|���F��/f_3���'�f*������o�n!��������ql.h�����`�B�ڛ|@����d���Y�a3���n m+��F�he�u|��
�L6�z�>>��k�.k4`oA�Ͷ�7C%����j�UUU
�`M�����@$e�����qE�(	* �i��H���'8�4`z�
>{�kT6�It^�K9��DX�u|6�Y����&K�1���w�Dj�s�b�o��e/�V4��!�_x���&��i���b�S�ф�9�ӣ��y��Z�\�(i�7b����>}�T�E���F���j���,�A˥7Ң�	{<a���\�+%G6Z"�W��d*^��g1��:{Px��$Y�l5�y([Tm�R��k+±#?���JD�l��Vt��Sh�,���*��*N�w!��+6�{i�݅ȦWN��a�v)��A��B�b*�gn@;��iB���9��WG�&	u��yƣ��0�
��ˎiF�Y�V�dx�5�W�Z􉵂b��Zm�Z6goX�j��p��2m@B1���;�����v��q�`�m����!�w�>a�#����A��.1�,�n�j��T?V/`y,�Ri�e��!�e���I`iQ��6�(���EP�m]&21���bf0=-`Q�d���&m���YO�4��&ֆ�}Z�d������x߯[MH�`����R'�j��M~ܱtV���4Y��g��i�
:;8\�ŏG�������6ՕY�cb�}J�9��^]76�k.|��Lu��/u�F?��6莊�,߇{Ԭ��e~�y'�'H��ҕ�rtF���{�ܙ~�����r�,�GRZ�{/N�����;K\�s&�i���xjt��>*��'�������Ψ���+FǼ��4L�	���L!	8.X8�(qϩB��%���`+�!�4��m�ڠc���u)HK|9����6E��2�E9bӃ�݅0�A�1w01�D֓,��e�6��!�q�0i�4�!��o�J���*�M'l��5$Шb�yy��X�)��c'ã���T���܈�}����!�Ud�t��<nB9�(� d�.u������[Տi�S�خ�S��#n7>Q�푦'���翩t��lT�m�4[��m�n}nf�NQM��f�Z�cC�#M�r�]R�*Bŋtp�zz�1�Sj��Y����c�EԚ0�j!�|G���}b������Fs�a�'�������SI�Ȟ,S0��E�ھ��*o��4�0��Q��\ʒ,~�§)@���1� Y<~X|�F��Q��v1V�F��E*\��� l40�TCK@��Ah(�k?B�]&O��%wj����0�ޖ�)Ij��ы���o����6��4��İ��9o��Nz�n���U=3�ں�U,��ߜb���Z"�Mf��l��#�Qk�=���h�L!)O~���{1�y��������tM!����Cs��-�c�J�X�HgA$?�M��\� !��u�X���m_V�	�L0�;"�aV]���ɢ+X7�q����w9����+Z;PC�X��m�d���1��O>����4��C��Mu�e��;,�г�+���W��.�}ꉿ�S*�Ҕ�{�a�/zΓ7�Ô�NJx�Yfٱ�s��1���t��e�5�I��y�L�]N-���B�=�TPS��tq�����"�(Hw����