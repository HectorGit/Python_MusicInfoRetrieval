BZh91AY&SY��oO �߀py���gߴ����P�띹��<ǒ5�UVR*~��G�2h    � "�P1     )�B�� � z�    E����)�dқ�!�6�ɦ ���z�D�&�x��S�*~���0C�4i��4�4*��ڈʫr���@!��������#��n�t�Z0���Q�
"���;XS��?�fQ�p���A�&(�$ǒ���I�si��?�^`���_B�^��˅qi�+���`���r"����k�7��&������Z1��ȭ&�ɭ.W+f�I ݊e���M�Q\0.�ı�(�L8<�&)�u�!#IǠ9B�����{ �>�hR��`����qynWV��,��=��/1ߥ@0�L ���all`$zFq9a�x-M4)�*�X!P �JrC����X�)��0�DD@q̓�!6�$z��a"Y�������5*�E�f=��N��T��U��E��
�M-��>��䐡	.4����	$?Cɵ:�F��U�/���
A�L�"�V���JJ��Ɔ!�͐�M
 ��d(&J(��%=L�p��,��eWw/K�4�jih�s����(.6yu���y�<�) ��R�#ȋ��~��ds��c@n��f�G�3��}�̽Ok/K�ё�C�Mn�S��+>��Q󁹴@rH2+�w��Z�GSĕ	yh��׼�r9 ]��{��P�8�s	��ima�K��b�M7���Jl|���C���^MM)WW>�цR�w�O�H��dì!J0��`(�Y[3�ųC�1WpbgX�$!$d!(�d����:��K{��m�����F��d��WZ}D�Ά��xx87>��y������d��A�R%�(��o
�Ě%nr5K	"io���
�Kxw:¤���oH¬���I����w��р�`F¬�5!!b4pZ�j�A�
2�qA0�!�\���z�:�#���-F���HY�F�K��XBD�@�G��D�u�G/=#A6��ց�z���:6���h;rz����4 ����Ϲ{�6� N �����e�z� ��/3p��R����/��������bY,�!�i�W&���Gm�48;���w�����m[��^�sŀ.�w��LO'�4��⁵�`�u�;B��cV��`����G���2M[����~.<Hh����{��|�:#�9!m�����<0Nx9I�.�p�!��ޞ