BZh91AY&SY��
  �߀Px���G߰?���@�8�:5��B=G�bf�Cj 444��4�4������h�    4J~�OP�=i���$0F�d�D�Ȃm*���j�OM=D� OD�W����$�<��J �e�6���a�;�G��?�U�ڣJ�\�W?y�Z�w�Ka��ӔyP�ō���u��eu�U�Gj�; �]�+��||}��/�7��ER~�%%#��5&�'!�Y���VT��e��"�ZF���4IPD���%y�Oe�Zp���F(�C�� XA$�a�Np����)';��ڊ�_�������zdt]��O'T��"������R��?g��͛�������P<B]�f9sZ�ٖ�g�+�f�Y���[�1a$�hd�Z����9񠈎�U/"��=���z'2m-ȄӔ��K/��:��q4��㠞���ԽB��,����q.�|���fV�K�l��hR	* �Ei�,S(���t����u���-)�U0�-�ͻM�X�9��h��j����D\B!�go)�3L��Ǻzf+nt jIT'k�&��&�+IF@߸�#Wl��"΁T��OmB�"H��b�Ֆ3�� ��xz�Ć�|�͝�CV�2*�C��im� b��Zɡ�1WF8d'��Q��#�xL���q�,��@���,�e����"3*�߆�^�մ}J�2�߫L� _�)�rE8P���
