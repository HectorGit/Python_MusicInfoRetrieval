BZh91AY&SY��� ߀Px���gߴ����Ps� c��d+�%	1&4S�m4)��zG��L�#OSi��JzI���@ d  h�BODQ�1M=@i�� �  昙2h�`��` ���D�#M&I�j6P<��d46��@��@�$I%`	@'����;
P�+c� ���;��I$+
3��{-<.7��,sٝi���   B   B ��ȗ�R����e���z�*)i��IN���/��2�md��uSOT����8DbpH���ݙ��<L��A�]œ�B�$��c@=/{kM�tۻb��ٙ�������ٚ.�n��^P �n@:H�����#wa�|Ps�'6�Ui^�2�؍���ip�[��Ēx�4�I�M�=rQl 9�"IqT�l�̺�@�$5��,���V]���K+E��,�!\6@F���$�U��Kwbm�V)���DJ���&">%�-����
I$�I)�Tі�fU��L�X�+۪�*��]��`D�.aC�K�2��P�L�y+��/��kn�s�6��5\�*ee���]��eyti�tߓ�r�A ��$J4��o?p��������x�| ��EW�xmgM�4&!��*&8��J��q	G���+Ǳ�ǜ@��%K�j]���x��Ɗ6w�ǭ�]����/7j��O��惮N������#GI��b�\�~�n�6־�B�* ��˗��/�=]�4=T8#Ũys�4�K�Q29�I�í�W��Y� �����UYǩ�&'N
�O:o�+7.�&UF4tK:�;eӢ�zՓ�N�8�Y�i���H�(�+�n��l0? (LM1�NeCpå[��ԙ�yU3�����N���S ��@�8�i���K�ytE8yȵ?u�g�3�q��;�2. GEE��m+��Ǚ(0�%�z|g�5���I�V�Y8��@�q ���i$J�Ԑ��Z���栲| �D���
�zK`$�8+(j��0e��'Xo��˘=ą��ƥ(��u��B0����'�Qgрcv��eC=U E�ڞ�NÆp��H�qa54l�5f���j�*�X(���ڻ�Ë9�N�q|����H�hɸ�R�!B�3_Y ���
cXF)n21���VD
���aI���B��F'	��U7$�3!?5,q��T�^��种]R5��(�J�S�rE8P����