BZh91AY&SYa�lg �_�px���o߰����`	_�׻) M��M��VPM�4OJy�z��6��������f����L�� &L   �� `�1 �&	�!��L���Sڔ=&�  �F��  9�#� �&���0F&"L��=T�I�OS�)�# �i��J�!j�@yA %$. $!(B��|�����4�$	�0Kރ�Ѷ�$�F
�H=%�%\B]���Q�q�eי-�����#�!A�f2%1�3�WxWy����ԩR�J�?��l{`�����q�ǓCy�M5�a��HQ�eS{)�3)��A,ɆP�L2-5	���]4"Sm�\B�L��V��-˶P��Ib���X���4aq�e/���C�rg";�n�k�X�vf���P��=�Ԟ�8 $pNԗ���Q�����L�M�R+��>�"�ɇ���J�$	ƦH�	P��]��O��ݦ�"��1���.	 LlE��|3^�V�#L�dF
NJ���H��Ѻ	$�"Z��"bt�kp�**�J�Z˰�&�d�2��1d�\wR�`�|^k��Clīx���(VԖu�$�y�ü��q�UH����)�:<��Ƶ�����$�2�Zb��օ��V�&�f�����Rv�[R��H�Uc�L�E�'Ʒ��ㅆ���Z8"
8�>�-�3�Ѷ�%����bm"�;��H��߀�VQS[ѧ8>ǽ��Κqơ0�N���q�w�pj���9;1�:;o]r
)8?%�9��AU�'gfN�1���Kr��N��5!1BL���
f,�*�ZL�����j�`���fd`�$@����H���CN�f�s����5F2H��|z�\�zy�X����s�Ծ��kH��Y�;G& �@�^䳘_&2!�mwV`�	����cf�0�B2�Z�-Qڲ��Q�͆�"��MQ�����_[1��]�ԏ��a՜̬�u�q�j�X��qsR	w'�	+��wB(��.5��݉$�K���tr�������F��W���0�x��b�]D�7��ɶ64�a���
;�ORӈ���|劄�%�	��^��*T��S�
�HXm�$��hc�L`�A �&FI%���Lc�,R�
*�J)P2��1*B`PA l<Y\�B�v��SMg��:�LhI6��<K�����ht�K<�5��]��$#��',���������̹K0XQ �� �pw��xɘe�~��1R@�͌ڍ������R24�$�0<ϻH�y�J�#�2��r_��!��.2���7�a�`��&�:׀V/;���ka��ؽ���P�u՚@ϒ��o}R��������d~���V;�f2KG�8I6�J�`^ ����`+�AG"TjI�������G�H�ơՙ� �$J
�@���ěD�FY��8��5�{ؑ}���7���WAS���������|���L B�@x�`��mD/ K`��nAB�(/ǆ��ay8$�Ug
��kM���qY#�KL��%� NV0&A�9��e�c�g3 ��v�I.i ]��Hj�z��;`�j���0H4�����P� ���tn��5!�	`8ҫ�T�
�\�.WF<�&b�Y%d��R��+Bn��KI���@�
����L�gA$x����YZOs@��L�MA�jjKj�փ4D�s6�$Q���rS�ѩ M��"�Z�l܍	 Y��>��iB�C�ma!�guV"�*���\��-�;+��60s�5�U��,�=cۦ�� WY���m�Vᶼ����� ��J�][�)Gˬ/�4�`&�9k�F ��=2�d�G0%����P2S�M�-�J�
�d�r(�'n�wWV�wWe�]�����8�>5�a!&X��rE8P�a�lg