BZh91AY&SY��~� �߀Px���gߴ����Pe�K�ֺa(���Q鲦h6�m5��4 5<��D����P�h  ��JPh � �   �12dф�14�&��	��x��d���m)�0�F���OQ➤��P"%D��
>����>E(?&*����<��RIh(ϣG��ZB_���ݬm�����w{�����y��M�5�0a��	�Z�b�Ή5k<8�v���Pa#B�8���w̝��Q�,�B
Y��J��xSL�g 8B�}"��l�4d*�1q6
��
�X�,h	yY�/U�����,u�kDh�]'bʄaZT���P�d1Q��1P�FUZ�HrsgpdVok��!2���!C0����K���>O8�I�O1H �liFナ�����:��5�q�)$��96�,i�ʩ��/C�SG"���=�@M)MI��s����{co_��J�-�=��=5>��ٰnL��ߣ?3�D	��w6�qL��&vMNƬ�;d�T��Q����
�TZ8G��ǘ��6kD�ڢH�v�����+��y?�9���#8K*3@�h���Ww��l��"cÚ����J{=<''
���Ja�]#&�l���8�I+���^jgհc�M��`Ò.n��g^�g��O���_?Vi� �A�H�C��_�Z��k(l�ad��/+���ǑCx�� �w�6g��u��*�����$:Og�0�o� [@9vji���ɓV�BqCb���A9��!�H������py�X)!�Cth�f�q,�ʸ���i�KQa�V@0�2��?���>�} �����JP~��ѿi%�/��ao;�q�XI�L� �@�IN۸3�#������|�n,l�#H3� ��ˆ��v[U$��\�F�'�<�l5�Q?�� ,���6�`2k:�U�Ϡ�v���J���00�/=^�|5HZ~^���HE���y�z*���f�My"cQ+Q@��h�rE8P���~�