BZh91AY&SY!-� �߀px���o߰����`	��u7�]{���Aϕmn�k�h�� @ �T���m'��1������(ȑD4       �{D��       ��EOЙ=C�!��2CF#ЁD�F�4&��i���F�1S �� �m)�l��mMM�h   *�8]�P%P�
,�G�9vU��Db�S)�$�����1J�'��BuB���p|/eU0�e��ŷ�q��Ӟ�����W�H����u�z�ɫ�t��"���mu��7z��]�{�ׯ�N,��s��:�~�>�,�6T��9������F�b��4x�"y�;��	fVe���e-Z�C£�C�����jnn�ǜ��̱�S)�C�tU��P�
R���ç�gA��ʸ�KT��SBq�j�@d�L#"4��DT0Ьa0�Ê����O:aC�i��� d��L��@�[)9�F�;��qN�'�� va�O���>#^,a33333 �����.�1���(Ƽ\��2HM��f�s��w�ަ;��Kq}�>�M�&�am���V�3T�d�4eɭ4���Uz�b����N��a�[��ؠ����U�P�r"e+93a2Fǵ]�ܵ�lP�EJé���U.�k����nQ�8��q;j˦�P2r�SDe0h�:P�K�*?\Tt���%t0��i*�1�e:pu�W����wKm��[ڲʆ�2!u7*�6�ΤCD̔?%�TR��f С�d�EXa5��X55�t�9����\��;P��+��L���
>����t�
�ͪxȊ��i8�QJ����i�� ���g'GZl�1��;_p�%��ih�U-#i����(�e�UEeU�McX�KP���VfF��%D�IJHK�Q�V�����b5E���JǬ�ئ&�jr��wв�ٸZ�I��K�J)̓�X�r�1 ˋ�'De����dC1�N%�S2'f�1����Ò�5�Cc��5�´n�DLZMMd5�X�e�|�';�7�8��i|���[�,���,,���V陷��t0��ᄕ�ޮ���.��tj�UUqW���s�*�N͏:8��۫-��I�3��e���}��|g���1UU�#Bx'G~D�����^������ؔ2�%)����n���1㩌�MՕeIL"��U@�uW�\,�eP�2UQPFn��C|�`Y�P�eZ)�ܫ�4!AH��%\�t��݇���g/�{,��H�!���'7w��Z]�%]}��Xx�H����p2O���nZ!5���4�϶G��[ھ/�^��s�-��y�V0�O���6�&%A�;OgR��q�/�5A6�T<��t��f�n����ސ�YS(c��ƫR�1#R__�/:iKW��m��1!�D�U\(p4Y���l:�'�42��� c툟t�:���k�"8E��Og	���Z��������J@S��gt ഢK�C&��z�;]�8�}SP��~�����
v�*0@���q�)�KE�er�H�kz�X���ʂ��(wFm�4���' �����,�\��kt;5��kz�ܘ�Rv
ܩ8�n���=f��$g�,`l*����"��6h����$T����=��H~�w�#3qHiow��]|��y��Rn ˒f���dcA�bI�\2���eD�C��W1���I\
�6��خ��+%r�bDU�Ĩ�4�ԓA�MB��o<ڥ�&.j��,��FH���mغ� ڳ"I M��@Kݽbb�=�燲��j8�.�.�+��L�w�3:dc����v�� ���!����A��5��e:F1����*�z�iKQ\�0�Q`�ۣ�w��\ۢ�� i��ڟ��M1����������Q�[�IE�q���uI����#q��eG��i.ihr�jh�Yq�jͤ��X�Υ���f������Y��#��'�ރ,�Ew=o���T���C�_�ף�nfGj,�%��ts�P�UXƀ����rE8P�!-�