BZh91AY&SYBF��  �_�Px���G߰?���@�DS��В$O)��&�&��fA��4�4�	M&�$��1<����y!�����`&F F&&	�bi�� �&&@     APf:	�DN�y�����fA���?~�@~�meJ,��ٍo[�<�Zn�^�nl�U���P�lQ�M�n���b���]���N�m\:��>nhE�Hs��L&Ύ�Q4 ��ކu�B��~���i���<�^I��1�2ޒI�i:CXڲ� �'sl�xB��B�0ͽ5�>� `��N��/�=��cV~�{	�;���5?}�gՓ��{��qտm3��8'<��$0�K�sY�`����]p�3�.�x;�\��k�ej��*��*OBm�qQ��m(6\�fD G��q�}�i��)��~�����8]13%��4ӽ�7��|d_H�)��h;�&�Zm�eK�XB[-�x�m|3���H,D��Vq��j Q)�
Rf`� =mx�3�Q�uw�)�$W4ogb댣+q2F�t�9inT���"�fGa�"d9��&$�8�ьl�&�5�,��j.FAeF�G������1�F�	u�bY�㷺��m�n��)i,wj�M�D�rhB���m���Bگ5�f�m�Z�9���9�P�׮���NUM$5J8����;�'^!e�n! �.KH	x?"1rE����X袊�u�4���*Sŉw�=#´_���"�(H!#ec�