BZh91AY&SY;�Ad _�Rxg������?���`�Ic��r�Ѡ 	!D�14��m��6��M	�?SDh4D����� h   �#!�4a0F�4b�20 JzJi4�� h �  �220CFi�F i�# ��A���L)��M$�j3Q���z�I�i��6�r ,�`�@M$�YRhGfHa��	"L��ҹL�M�2iɏ��*�޳�oE<K�?|�TY�{:�X譑���t�-ImF���;͔�8B�f�0:���?(F�X����� ��&0ͯN��g�#�\�=d�W���]m�g�0�[
�_��Ղ�S�]�O�����㍜�X����QvQ0���H��\]Z�6o��O�/��(YE�gSIB���	@dm�������*̴�X�np�N�~#;�.�B��T��;ϙ��VyUr����[Fcl�kG���0i�7>z���x�4`.��c&��r�FY�<�Ĺ�V�U���e��r�,����qu�p�|��2�<��9�ؗr�k=���#Q#�Oѣj�yv��Y2���!����)���u����������F���=�auB��J��R��@�R6$�b�V�P�J�-NV��ac0R�4`/Il��Y�`qX�C|��Z9.3	�q�9�5����#)B�E��j��\5���i���0�zq�dŠ,��wy�����N�0眇�n�0fA"%��0-j��R��Ҍ���#P|pm�bU��e6B�{@�V����JKaNɓW$�V1�fa�Ao�a�DlDTMB#�9UZ�ֆ�ئ�(C-D.U�4F��!�h p5�5Q��	
�k9��p��������X��:�s������˫�&�FK	��~�C���$���6��+�ZN9�-��)K(p]�d6]MJ��c�� ��u���9~n�7�QXL���䴖��[�Z��a2`.����w2�^��i��	t'L�N�
5��a�څ�>�qK2�9ye�(�~��Y���؍�C$
E�×�g�'�jH֏K7��A�)���$t�S���`�`�7)�)a�Ab��=̂aB��2��S��,�I$��|.��@�.vH��%D��^�r2��!x	�D��3���"��B�8�cB��k�%��MeR��-@����lV>��ԓH��C�+.K�����`��  Z�����V��I='�3+X�O[	ç̰
H㶂Jǡ-oעF�uX��	"G0��$#� 2;k�+�t0�T�FfSG��k��܊P������IT7ƙ�*�q�h�O��9!��B��q.������cL�Ƅ@@G6e�;w��*�	�e�� W�������X4�P��$~Ǭ�*x0Jm��
i��� i&-��
��&d3"lsL�F�(@�!�����8g���bT>M慆�*��c
����7� δ4j	�AkX;�D1��@�*��4��H�"	���m6���p���	>�U���L��Y�&0%�J4����?v~҆I��LMa dw�7�v�ަmh����]K��J M�K�]�3��!$A��c�@�6l�N��qI�%4$�;Ť���9Ci���
&�������TS{���*N�Ra2Q�Ҵ���f�hoQSy��p�-)R��C"��bT�sD�7G���E�U�&0���A��CF�@�[����Μ���R��Y8b$b�6p"k
{��X�:����1y���cB��s���L��=�ϸ9�� �@���z;[V�K3�7"�E�1�\8L-�W6��ugY�y�x�'�������2�`Yb�H��rE8P�;�Ad