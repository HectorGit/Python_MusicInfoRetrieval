BZh91AY&SY(� � �߀py��O߰?���`zۡ� �J �Q��A��M  Ѧ@  hjJ�   �LM��&MLL`��HH�M&��&�d	�����d`M2�&MLL`��E AM1���� �Q� �M=%0nI
`�O��VbǏ����a��}�dB���H=��ZZK��r8�8����v��}��ul�OI�Y��AHdD  z�f��"p�"��*X�b��1�Am�5vy3����!-��:�ed�ܳ�kYe�52	)n������}w��I�9Kgb�ၛ�w1G������P2qڜ�Z�.4��VS����������]�xx�����@ o7D$f*9�n\r�8`����8$c ��L�U�*�ց�U��T��br�\��H�o'2�R��(6�-i� ��1�'Q�b���Rr�RH��#e��c�ý�o/�XR�.G`����s�tBt
?X!� !jvb(4)#:l��Ju`%2"�m� ���M:�"mQ�J�E5��Dp���J�X�ddE8@E�<q���Q`��7�z��Bقz-T�y��� ��5Ze|6���I,��­���5�X���8)�<��`66#YyŽ)U�� �ab�C���XT�Cl�)+���(ܝy�������$�B�F�,���/�I��m�����?5�\��u�K�(B��x�!E����|��`������*-�#y�Q)`Fl�c#f��p���E�X������XC��#�'G7;�a�Z
���j�/̼��i�2�z0�o"�X$���'lsXm����i�aՋ#y�f�Y����x:NA��?�6�`Ē�9��x!1.�>d���&�̒�H%y*�.��R�0X*�a����v��h��cfa%7#�`�$Ca�g�ef*V�U*DR�r���1��d�
(-Z�Mo���,�r=:��/)�8��lz�:����G�Ժ������թ�e��a�.S�젡e�4��8�������}oă � U�9;�w�F�;���0���iv�*�>{c#�A	�ȴ���C5��?>�`�Y��$΋�e��n��V�3�<����H	��AI ���� ��Э��"��rT�C���X&T�`��4&�F�[��X�?#�^01�i`��9�66=g�;2`  /(l&� �x�<��03T�� ��^����pҩMF��,t{�lƂX�^u�zp�F�>�^W�;�=h��%P�{C�
��s'f������ȄRa9���aLT	�</3�͋�����I,����6��6
Zd�"&��#���\�m��_S�Pq��t��|��e��m8D��s��Fc��v+�Hv�B��x@����V$y��������&F�D~b8��� �T�аL�}%�5l_�z�#9ӨR.���I�".�	�eN�Et�,j��{�<1��iA>��"F�9dC�&�AD�<y�}��؏i��13^�"�3��c�hjg?�w$S�	�`	p