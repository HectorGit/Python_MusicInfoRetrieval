BZh91AY&SY���� ߀Px��G߰?���@�� G0 L� L&	�0`��S�@h�    s ɀ�`�C F 
�&��К1M��&����4�4~���]��B�^�DR"�G��RJa�syID#��[R#��g��ID�iVkV�#���>m	JK꺎�pV��Ǡ��_$W&zM0������Kp�wT�9R�Ef"Q���m�rK$�k�2���PX1)Ha[��6��Y(��I	W8����y%J.\�s�b�w]��ʨ�U���bI@iF(JB�D��d�Wu�2���h�iy��b�o�k���(\���U[�x0�s����>��wtw#SGs�F���.�.y�9�*�w�D`�"����b.�oͺj�KbZ_e"[[��M��]���a��y(�h̹�B'�2;��ã�n���D��&��7�W0mԊ��U��m٥�C����t��#�o�9�_�oY�-�����rF���l�-{������(�bR���tFE_~Fj��NJ%0�F�O��Qe(Х�j�ՠ�pU���:����d=/�8�*P���[J:��a2���\�lWŌ;)F�p�Z�|}X/S�J�K�+K��Lhe�N��ʸ��jT�FN��7��Άb��!��V���&P�1�0�d{�(��(�7���rE8P�����